<svg width="617" height="173" viewBox="0 0 617 173" fill="none" xmlns="http://www.w3.org/2000/svg">
<path d="M194.165 122H214.405V84.5835C214.405 83.5825 214.265 82.3213 213.984 80.7998C213.704 79.2383 213.544 78.1772 213.504 77.6167H214.285C214.485 78.2173 214.865 79.2783 215.426 80.7998C215.986 82.2812 216.527 83.5625 217.047 84.6436L242.812 122H263.413L289.058 84.5835C289.538 83.5425 290.039 82.4014 290.559 81.1602C291.12 79.9189 291.56 78.7378 291.88 77.6167H292.661C292.541 78.6577 292.361 79.8188 292.121 81.1001C291.92 82.3813 291.82 83.5625 291.82 84.6436V122H312.721V57.0166H282.691L256.626 93.1719C256.105 94.2529 255.585 95.2939 255.064 96.2949C254.584 97.2559 254.124 98.3369 253.683 99.5381H253.263C252.822 98.3369 252.362 97.2559 251.881 96.2949C251.401 95.2939 250.88 94.2529 250.32 93.1719L224.134 57.0166H194.165V122ZM323.051 90.7695C323.051 101.66 326.614 109.708 333.741 114.913C340.908 120.118 350.778 122.721 363.35 122.721C375.642 122.721 385.312 120.118 392.358 114.913C399.445 109.708 402.989 101.66 402.989 90.7695V57.0166H381.788V93.7725C381.788 99.0176 380.106 102.741 376.743 104.943C373.38 107.105 368.815 108.187 363.05 108.187C357.124 108.187 352.5 107.105 349.176 104.943C345.893 102.741 344.251 99.0176 344.251 93.7725V57.0166H323.051V90.7695ZM410.856 103.682C410.856 110.048 414.56 114.813 421.967 117.976C429.415 121.139 438.964 122.721 450.615 122.721C462.307 122.721 471.696 120.939 478.783 117.375C485.91 113.812 489.473 108.767 489.473 102.241C489.473 96.5952 487.271 92.0708 482.867 88.6675C478.462 85.2241 470.214 82.3613 458.123 80.0791C448.033 78.4375 441.186 77.3164 437.583 76.7158C433.979 76.0752 432.177 75.4746 432.177 74.9141C432.177 73.5127 433.599 72.4917 436.441 71.8511C439.284 71.1704 443.789 70.8301 449.955 70.8301C455.92 70.8301 460.445 71.2905 463.528 72.2114C466.651 73.0923 468.212 74.4136 468.212 76.1753V78.2173H487.191V74.4937C487.191 69.2485 483.728 64.9243 476.801 61.521C469.914 58.0776 460.845 56.356 449.594 56.356C438.223 56.356 429.174 58.0776 422.448 61.521C415.721 64.9243 412.358 69.729 412.358 75.9351C412.358 81.1802 414.62 85.5845 419.145 89.1479C423.709 92.7114 432.197 95.6943 444.609 98.0967C455.14 99.8984 461.946 101.08 465.029 101.64C468.152 102.161 469.714 103.021 469.714 104.223C469.714 105.664 468.032 106.785 464.669 107.586C461.346 108.347 456.581 108.727 450.375 108.727C443.969 108.727 438.984 108.167 435.42 107.045C431.857 105.924 430.095 104.183 430.135 101.82V98.8774H410.856V103.682ZM497.761 122H519.322V57.0166H497.761V122ZM528.331 89.3281C528.331 101.5 532.355 110.188 540.403 115.394C548.491 120.559 559.381 123.141 573.075 123.141C586.007 123.141 595.997 121.379 603.044 117.856C610.131 114.333 613.714 109.107 613.794 102.181V95.8145H593.735V101.34C593.935 103.021 592.494 104.683 589.411 106.325C586.368 107.926 581.143 108.727 573.735 108.727C566.809 108.727 561.283 107.746 557.159 105.784C553.035 103.782 550.973 100.359 550.973 95.5142V83.5024C550.973 80.8999 552.975 78.0972 556.979 75.0942C560.983 72.0513 566.508 70.5298 573.555 70.5298C579.921 70.5298 584.546 71.3706 587.429 73.0522C590.352 74.6938 592.394 75.7749 593.555 76.2954L593.735 83.5024H613.794L613.674 78.2173C611.592 70.2896 607.508 64.584 601.422 61.1006C595.376 57.5771 585.947 55.8154 573.135 55.8154C559.922 55.8154 549.151 58.3579 540.823 63.4429C532.495 68.4878 528.331 77.2363 528.331 89.6885V89.3281Z" fill="white"/>
<path d="M153.5 75.2417C162.167 80.2454 162.167 92.7546 153.5 97.7583L62.75 150.153C54.0833 155.157 43.25 148.902 43.25 138.895V34.1055C43.25 24.0981 54.0833 17.8434 62.75 22.8471L153.5 75.2417Z" fill="white"/>
</svg>